module sqrt(a,out);
input logic a;
output logic out;




endmodule