

module divider (a,b,out);

    
endmodule
