// module multiplication_normaliser(in_e, in_m, out_e, out_m);
// input  logic [7:0] in_e;
// input  logic [47:0] in_m; // as the product of two 24 bit no's is 48 bit wide
// output  logic [7:0] out_e;
// output  logic [47:0] out_m;


// always@(*) begin
    

//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end
//     if(in_m[47:0]==48'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001) begin
//         out_m=in_m<<47;
//         out_e=in_e-47;
//     end

// end






// endmodule

module multiplication_normaliser(in_e, in_m, out_e, out_m);
  input  logic [7:0] in_e;
  input  logic [47:0] in_m; // as the product of two 24 bit no's is 48 bit wide
  output  logic [7:0] out_e;
  output  logic [47:0] out_m;

  genvar i;

  always @(*) begin
    if (in_m[47:0] == 48'b0) begin
      out_m = in_m << 47;
      out_e = in_e - 47;
    end else begin
      out_m = in_m;
      out_e = in_e;
    end

    for (i = 0; i < 48; i = i + 1) begin
      if (in_m[i] == 1'b1) begin
        out_m = in_m << (47 - i);
        out_e = in_e - i;
        break;
      end
    end
  end
endmodule
